module porta_e(A, B, S);

    input A, B;
    output S;

    assign S = A & B;

endmodule